[aimspice]
[description]
281
Redresor cu filtru

D1 1 2 DiodaS
D2 0 1 DiodaS
D3 0 3 DiodaS
D4 3 2 DiodaS
.model DiodaS D tt=1e-9

C1 2 0 1m
rl 5 0 100
r1 2 4 220

dz 0 4 zener
.model zener D bv = 6.8

q1 2 4 5 transistor
.model transistor npn tr = 1e-9 tf = 1e-9

vin 1 3 sin(0 10 50 0 0)


[tran]
1e-9
60e-3
X
X
0
[ana]
4 1
0
1 1
1 1 -3.41661E-22 6
1
v(5)
[end]
