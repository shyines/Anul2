[aimspice]
[description]
228
Nand:
.model nand nmos vto=2.5
M3 vdd vgg vout vout nand l=25u w=10u
M2 vout a x x nand l=1u w=10u
M1 x b 0 0 nand l=1u w=10u
va a 0 dc 0 pulse(0 5 0 1e-10 1e-10 1e-9 2e-9)
vb b 0 dc 5
VDD vdd 0 dc 5
VGG vgg 0 dc 7.5


[dc]
1
va
0
5
0.1
[tran]
1e-9
6e-3
X
X
0
[ana]
1 1
0
1 1
1 1 -1 6
3
v(a)
v(b)
v(vout)
[end]
