[aimspice]
[description]
373
Redresor cu filtru
D1 1 2 Dioda
D2 3 2 Dioda
D3 0 3 Dioda
D4 0 1 Dioda
.Model Dioda D
R 2 0 100
C 2 0 3m
Vin 1 3 sin(0 10 50 0 0)
!*Condensatorul inmagazineaza energie cand tensiunea furnizata de redresor e mai mare decat cea dintre armaturile sale
!*Condensatorul debiteaza energie cand tensiunea furnizata de redresor e mai mica decat cea dintre armaturile sale
[tran]
1e-8
60e-3
X
X
0
[ana]
4 1
0
1 1
1 1 -2 10
3
v(1)
v(2)
v(3)
[end]
